module audio_buffer
 ( input rx_data, rx_lrclk, rx_sclk, rx_lock,
   output tx_data, tx_lrclk, input tx_sclk,
   output almost_full, almost_empty, is_full, is_empty,
   output reg overflow, underflow
 );
 
 reg [6:0] rx_byte;
 reg [4:0] rx_cnt;
 reg [5:0] tx_cnt;
 reg rx_lrclk_1;
 reg [8:0] m_byte;
 reg [7:0] tx_byte;
 reg tx_lr;
 
  initial
  begin
	  rx_lrclk_1 = 0;
	  rx_cnt = 0;
	  tx_cnt = 0;
	  rx_byte = 0;
	  tx_byte = 0;
	  m_byte = 0;
	  tx_lr = 0;
	  overflow = 0;
	  underflow = 0;
  end
	  
 // de-serialyze into stream of bytes
 // assume 'left justified' input format:
 // first data bit comes together with the first '1' state of the lrclk.
 // data and lrclk change at falling edge of sclk, and are meant to be
 // stable and clocked-in at the posedge of sclk
 
 wire       fifo_d_en = (rx_cnt[2:0] == 3'h7) && (rx_cnt[4:3] != 2'h3);
 
 always @(posedge rx_sclk)
 begin
	rx_lrclk_1 <= rx_lrclk; // remember previous value
	if (!rx_lock || (rx_lrclk && !rx_lrclk_1)) // start with new incoming sample
		rx_cnt <= 1; // counter contains the number data bits sampled in the shiftreg
	else
		rx_cnt <= rx_cnt + 1;
	// shift-in new incoming data bit
	rx_byte <= {rx_byte[5:0], rx_data};
		
	// copy-out filled-up byte: first 3 bytes of each 4-byte sample
	//if (rx_cnt[2:0] == 3'h7 && (rx_cnt[4:3] != 2'h3))
	//begin
	//	m_byte <= {rx_lrclk, rx_byte, rx_data};
	//	rx_flag <= !rx_flag;    // toggle receiver flag, assume buffer was empty
	//	if (rx_flag != tx_flag) // rx_flag==tx_flag indicates empty. A full mbyte got overwritten!!
	//		overflow <= !overflow; // toggle value to indicate overflow
	//end
	if (fifo_d_en && is_full)
    begin
		overflow <= !overflow; // toggle value to indicate overflow
    end
 end
 
 wire [8:0] fifo_d    = {rx_lrclk, rx_byte, rx_data};
 wire       fifo_d_ck = rx_sclk;
 wire [8:0] fifo_q ;
 wire       want_sample = (tx_cnt[2:0] == 0) && (tx_cnt[4:3] != 2'h3);
 wire       fifo_q_en = want_sample && !is_empty && (tx_cnt[5] == fifo_q[8]);
 wire       fifo_q_ck = !tx_sclk;
   
  // mbyte async buffer control:
  // it contains a value if rx_flag != tx_flag, otherwise it is empty
	
  // on transmit side, outbound data and lrclk must change at tx_sclk negedge
  always @(negedge tx_sclk)
  begin
	tx_cnt <= tx_cnt + 1;
	  
	if (want_sample) // first 3 bytes of every (4-byte) L/R word
	begin // every 8th cycle of bit counter we can pull a next byte from the audio buffer
		if (fifo_q_en)
			{tx_lr,tx_byte} <= fifo_q;
		else
	    begin // insert silence on audio out
		    underflow <= !underflow; // toggle value to indicate underflow
		    {tx_lr,tx_byte} <= {tx_cnt[5], 8'h0};	
		end
	end
	else // shift out serial audio data from byte buffer, also 0s for 4th byte
		tx_byte <= {tx_byte[6:0],1'h0};
  end
  
  assign tx_lrclk = tx_lr;
  assign tx_data = tx_byte[7];
  
  
 /* Verilog module instantiation template generated by SCUBA Diamond (64-bit) 3.3.0.109 */
/* Module Version: 5.7 */
/* Fri May 01 00:03:05 2015 */
/* parameterized module instance */
Ipexpr_fifo ipfifo (.Data(fifo_d), .WrClock(fifo_d_ck), .RdClock(fifo_q_ck), .WrEn(fifo_d_en), .RdEn(fifo_q_en), 
    .Reset( 1'h0), .RPReset( 1'h0), .Q(fifo_q), .Empty( is_empty), .Full( is_full), .AlmostEmpty( almost_empty), 
    .AlmostFull( almost_full));
	
// TODO: check and repair for the clockdomain crossings of the use of the (alomst-)empty/full signals.
 endmodule